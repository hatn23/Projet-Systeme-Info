----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:47:43 05/02/2020 
-- Design Name: 
-- Module Name:    MemoireInstruction - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MemoireInstruction is
    Port ( ADDR : in  STD_LOGIC_VECTOR (7 downto 0);
           CLK : in  STD_LOGIC;
           OUTPUT : out  STD_LOGIC_VECTOR (31 downto 0));
end MemoireInstruction;

architecture Behavioral of MemoireInstruction is
type table is array (0 to 15) of STD_LOGIC_VECTOR(7 downto 0);
signal donnee: table ;
begin
	process
	begin
		wait until CLK'event and CLK='1';
			OUTPUT<= donnee(to_integer(unsigned(ADDR)));
	end process;

end Behavioral;

